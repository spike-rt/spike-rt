/*
 * SPDX-License-Identifier: MIT
 *
 * Copyright (c) 2023 Embedded and Real-Time Systems Laboratory,
 *            Graduate School of Information Science, Nagoya Univ., JAPAN
 */

/*
 *  Pybricks USB用SIOドライバ
 */

[singleton]
celltype tSIOAsyncPortPybricksUSB {
  entry   sSIOAsyncPort eSIOPort;
  entry   sSIOAsyncCBR  eSIOCBR;
  [optional] call    sSIOAsyncCBR  cSIOCBR;
};


/*
 *  シリアルインタフェースドライバのプロトタイプ
 */
[prototype]
cell tSIOAsyncPortPybricksUSB SIOAsyncPortPybricksUSB1 {
};
